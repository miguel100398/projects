`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:03:20 05/09/2017 
// Design Name: 
// Module Name:    PC 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module InstructionMemory(
    input [31:0] Address,
    output [31:0] Word
    );
	
	/*
	 ROM_1 r1(
	 .a(Address[5:0]),
	 .spo(Word)
	 );
	 */
	 
	 
	 
	 
	 
	 ROM_SAD r1(
	 .a(Address[6:0]),
	 .spo(Word)
	 );
	 
	 
	 
	/*
	 ROM_3 r1(
	 .a(Address[5:0]),
	 .spo(Word)
	 );
	 */
	 
	 


endmodule
