module SAD (
input clk,
		rst,
		go,
input [7:0] A [15:0],
input [7:0] B [15:0],
output [7:0] AB_addr,
output [31:0] sad
);

logic i_lt_16;
logic Ab_rd;
logic i_inc;
logic i_clr;
logic sum_ld;
logic sum_clr;
logic sad_reg_ld;
logic sad_reg_clr;

logic [7:0] i;
logic [31:0] sum;
logic [31:0] sum_abs;
logic [31:0] sad_reg;
logic [31:0] subs [15:0];
logic [31:0] abs [15:0];

FSM fsm1 (
.go(~go),
.i_lt_16(i_lt_16),
.rst(~rst),
.clk(clk),
.AB_rd(Ab_rd),
.i_inc(i_inc),
.i_clr(i_clr),
.sum_ld(sum_ld),
.sum_clr(sum_clr),
.sad_reg_ld(sad_reg_ld),
.sad_reg_clr(sad_reg_clr)
);

//////////////////// i /////////////////////////////////////////////////////////////////////////
always_ff @ (posedge clk) begin
	if (i_clr) 
		i = 0;
	else if (i_inc)
		i = i + 1;
	else
		i = i;
end
/////////////////////////////////////////////////////////////////////////////////////////////////

/////////////////////comparador/////////////////////////////////////////////////////////////////
always_ff @ (posedge clk) begin
	if (i<16)
		i_lt_16= 1;
	else
		i_lt_16 = 0;
end
///////////////////////////////////////////////////////////////////////////////////////////////

/////////////////////SUM///////////////////////////////////////////////////////////////////////
always_ff @ (posedge clk) begin
	if (sum_clr)
		sum = 0;
	else if (sum_ld)
		sum = sum + sum_abs;
	else
		sum = sum;
end
///////////////////////////////////////////////////////////////////////////////////////////////

//////////////////sad_reg/////////////////////////////////////////////////////////////////////
always_ff @ (posedge clk) begin
	if (sad_reg_clr)
		sad_reg = 0;
	else if (sad_reg_ld)
		sad_reg = sum;
	else
		sad_reg = sad_reg;
end
/////////////////////////////////////////////////////////////////////////////////////////////

///////////////////////////Restadores///////////////////////////////////////////////////////
integer p;
always_comb begin
	for (p = 0; p < 16; p = p + 1) begin
		if (~rst)
			subs [p] = 0;
		else
			subs [p] = A[p] - B[p];
	end
end
////////////////////////////////////////////////////////////////////////////////////////////

///////////////////////////Absolutes////////////////////////////////////////////////////////
integer q;
always_comb begin
	for (q = 0; q < 16; q = q +1) begin
		if (~rst)
			abs[q] = 0;
		else if (subs [q] [31] == 0 )
			abs[q] = subs [q];
		else abs[q] = ~subs[q] +1;
	end
end
////////////////////////////////////////////////////////////////////////////////////////////

//////////////////////////Sum_abs/////////////////////////////////////////////////////////
assign sum_abs = abs[0] + abs [1] + abs[2] + abs[3] + abs[4] + abs[5] + abs[6] + abs[7] + abs[8] +
abs[9] + abs[10] + abs[11] + abs[12] + abs[13] + abs[14] + abs[15];
////////////////////////////////////////////////////////////////////////////////////////////


assign AB_addr = i;
assign sad = sad_reg;

endmodule 